//    This is a component of pluto_step_spi, a stepper driver for linuxcnc over SPI.
//    based on the main.v from Jeff Epler <jepler@unpythonic.net>
//    Copyright 2013 by Matsche <matsche@play-pla.net>
//
//    This program is free software; you can redistribute it and/or modify
//    it under the terms of the GNU General Public License as published by
//    the Free Software Foundation; either version 2 of the License, or
//    (at your option) any later version.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program; if not, write to the Free Software
//    Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA
//**********************************************************************
//`define USE_SERVO
// Open-Drain buffer
//`define OD
`ifdef OD
module OC_Buff(in, out);
input in;
output out;
assign out = in ? 1'bz : 1'b0;
endmodule
`endif
//all = 31
//uni = 14 
// in = 5  + rpm =1
//out = 10 + pwm/rc=1
module spi_main(clk, SCK, MOSI, MISO, SSEL, LED, dout, din, step, dir, pout, rin);
parameter W=10;
parameter F=11;//velocity width
parameter T=5;//time width *1600ns
parameter I=16;//pins input
parameter O=16;//pins output
parameter INV_PWM=0;//invert pwm
input clk;

input SCK, SSEL, MOSI;
output MISO;
output LED;
input [I-1:0] din;
input rin;//rpm in

reg Spolarity;
reg [3:0] Dpolarity;

reg[O-1:0] real_dout; output [O-1:0] dout = /*do_tristate ? {O-1{1'bZ}} :*/ real_dout; 
wire[3:0] real_step; output [3:0] step = /*do_tristate ? 4'b0 :*/ real_step ^ {4{Spolarity}};
wire[3:0] real_dir; output [3:0] dir = /*do_tristate ? 4'b0 :*/ real_dir ^ Dpolarity;
wire real_pout; output pout = /*do_tristate ? 1'b0 :*/ (INV_PWM)?~real_pout:real_pout;

`ifdef OD
OC_Buff ocout[O-1:0](real_dout, dout);
OC_Buff ocstep[3:0](real_step ^ {4{Spolarity}}, step);
OC_Buff ocdir[3:0](real_dir, dir);
`endif

wire [W+F-1:0] pos0, pos1, pos2, pos3;
reg  [F:0]     vel0, vel1, vel2, vel3;
reg [T-1:0] dirtime, steptime;
reg [1:0] tap;
reg [7:0] in_pwm = 8'd0;
wire [15:0] rpm;

reg [10:0] div2048;
wire stepcnt = ~|(div2048[5:0]);
wire in_clk=stepcnt;//&div2048;

always @(posedge clk) begin
    div2048 <= div2048 + 1'd1;
end

wire do_enable_wdt, do_tristate;
wdt w(clk, do_enable_wdt, in_clk, do_tristate);
`ifdef USE_SERVO
rcservo s(in_pwm, in_clk, real_pout);
`else
pwm p(in_pwm, in_clk, real_pout);
`endif
rpm r(rin, &div2048[8:0], rpm);
stepgen #(W,F,T) s0(clk, stepcnt, pos0, vel0, dirtime, steptime, real_step[0], real_dir[0], tap);
stepgen #(W,F,T) s1(clk, stepcnt, pos1, vel1, dirtime, steptime, real_step[1], real_dir[1], tap);
stepgen #(W,F,T) s2(clk, stepcnt, pos2, vel2, dirtime, steptime, real_step[2], real_dir[2], tap);
stepgen #(W,F,T) s3(clk, stepcnt, pos3, vel3, dirtime, steptime, real_step[3], real_dir[3], tap);

//**********************************************************************
// SPI zeugs
// synchronizing the handshakes
//
reg [2:0] SCKr;
always @(posedge clk) SCKr <= {SCKr[1:0], SCK};
wire SCK_risingedge = (SCKr[2:1]==2'b01);  // now we can detect SCK rising edges
wire SCK_fallingedge = (SCKr[2:1]==2'b10);  // and falling edges
//wire SCK_high = SCKr[1];  // SCK is high

// same thing for SSEL
reg [2:0] SSELr;
always @(posedge clk) SSELr <= {SSELr[1:0], SSEL};
wire SSEL_active = ~SSELr[1];  // SSEL is active low
wire SSEL_startmessage = (SSELr[2:1]==2'b10);  // message starts at falling edge
//wire SSEL_endmessage = (SSELr[2:1]==2'b01);  // message stops at rising edge

wire MOSI_data = MOSI;

// we handle SPI in 8-bits format, so we need a 3 bits counter to count the bits as they come in
reg [2:0] bitcnt;
reg byte_received;  // high when 8 bit has been received
reg [4:0] spibytecnt;
reg [7:0] data_recvd;
reg [7:0] data_sent;
reg [7:0] data_outbuf;

always @(posedge clk) begin
	if(SSEL_startmessage) begin
		//data_sent <= data_outbuf;
		bitcnt <= 3'b000;
		spibytecnt <= 5'b00000;
	end
	if(SSEL_active) begin
		if(SCK_risingedge) begin
			data_recvd <= {data_recvd[6:0], MOSI_data};
			bitcnt <= bitcnt + 3'b001;
			if(bitcnt==3'b000)
				data_sent <= data_outbuf;
		end
		else if(SCK_fallingedge) begin
			data_sent <= {data_sent[6:0], 1'b0};
			if(bitcnt==3'b000) begin
				spibytecnt <= spibytecnt + 5'b00001;
			end
		end
		byte_received <= SCK_risingedge && (bitcnt==3'b111);
	end
end
assign MISO = data_sent[7];  // send MSB first
// we assume that there is only one slave on the SPI bus
// so we don't bother with a tri-state buffer for MISO
// otherwise we would need to tri-state MISO when SSEL is inactive

reg [7:0] data_inbuf;
always @(posedge clk) begin
	if(SSEL_active) begin
		//------------------------------------------------- word 0
		if(spibytecnt == 5'b00000) begin	// 0
			data_outbuf <= pos0[7:0];
			if(byte_received)
				data_inbuf <= data_recvd;	//vel0[7:0] 
		end
		else if(spibytecnt == 5'b00001) begin	// 1
			data_outbuf <= pos0[15:8];
			if(byte_received)
				vel0 <= {data_recvd[F-8:0],data_inbuf};	//vel0
		end
		else if(spibytecnt == 5'b00010) begin	// 2
			data_outbuf <= pos0[W+F-1:16];
			if(byte_received)
				data_inbuf <= data_recvd;	//vel1[7:0]
		end
		else if(spibytecnt == 5'b00011) begin	// 3
			data_outbuf <= 8'b0;
			if(byte_received)
				vel1 <= {data_recvd[F-8:0],data_inbuf};	//vel1
		end
		//------------------------------------------------- word 1
		else if(spibytecnt == 5'b00100) begin	// 4
			data_outbuf <= pos1[7:0];
			if(byte_received)
				data_inbuf <= data_recvd;	//vel2[7:0]
		end
		else if(spibytecnt == 5'b00101) begin	// 5
			data_outbuf <= pos1[15:8];
			if(byte_received)
				vel2 <= {data_recvd[F-8:0],data_inbuf};	//vel2
		end
		else if(spibytecnt == 5'b00110) begin	// 6
			data_outbuf <= pos1[W+F-1:16];
			if(byte_received)
				data_inbuf <= data_recvd;	//vel3[7:0]
		end
		else if(spibytecnt == 5'b00111) begin	// 7
			data_outbuf <= 8'b0;
			if(byte_received)
				vel3 <= {data_recvd[F-8:0],data_inbuf};	//vel3
		end
		//------------------------------------------------- word 2
		else if(spibytecnt == 5'b01000)  begin	// 8
			data_outbuf <= pos2[7:0];
			if(byte_received)
				data_inbuf <= data_recvd;	//real_dout[7:0]
			end
		else if(spibytecnt == 5'b01001) begin	// 9
			data_outbuf <= pos2[15:8];
			if(byte_received) begin
				real_dout <= {data_recvd[O-8-1:0], data_inbuf};	//real_dout
			end
		end
		
		else if(spibytecnt == 5'b01010) begin	// 10
			data_outbuf <= pos2[W+F-1:16];
			if(byte_received)
				data_inbuf <= data_recvd;
		end
		else if(spibytecnt == 5'b01011) begin	// 11
			data_outbuf <= 8'b0;
			if(byte_received) begin
				tap <= data_recvd[7:6];
				steptime <= data_recvd[T-1:0];
				Spolarity <= data_inbuf[7];
				dirtime <= data_inbuf[T-1:0];
			end
		end
		
		//------------------------------------------------- word 3
		else if(spibytecnt == 5'b01100) begin // 12
			data_outbuf <= pos3[7:0];
			if(byte_received) begin
				in_pwm <= data_recvd;
			end
		end
		else if(spibytecnt == 5'b01101) begin //13
			data_outbuf <= pos3[15:8];
			if(byte_received) begin
				Dpolarity <= data_recvd[3:0];
			end
		end
		else if(spibytecnt == 5'b01110) data_outbuf <= pos3[W+F-1:16];//14
		else if(spibytecnt == 5'b01111) data_outbuf <= 8'b0;//15
		//------------------------------------------------- word 4
		else if(spibytecnt == 5'b10000) data_outbuf <= din[7:0];//15
		else if(spibytecnt == 5'b10001) data_outbuf <= din[I-1:8];//I-1:8];//17
		else if(spibytecnt == 5'b10010) data_outbuf <= rpm[7:0];//8'b0;//18
		else if(spibytecnt == 5'b10011) data_outbuf <= rpm[15:8];//8'b0;//19
		else data_outbuf <= spibytecnt;//20
	end
end
//assign LED = do_tristate ? 1'bZ : (real_step[0] ^ real_dir[0]);
assign do_enable_wdt = data_recvd[6] & (spibytecnt == 5'b01001) & byte_received;
assign LED = in_clk;

endmodule
